typedef uvm_sequencer#(intr_tx) intr_sqr;