typedef uvm_sequencer#(intr_tx) mem_sqr;